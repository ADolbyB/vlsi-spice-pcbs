** Profile: "SCHEMATIC1-optest1"  [ C:\Users\JB\Desktop\Code\PSpice\homework1-pspicefiles\schematic1\optest1.sim ] 

** Creating circuit file "optest1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_DATA\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.3ms 0 1us 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
